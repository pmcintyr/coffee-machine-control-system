architecture rtl of bin_to_bcd is
    --It is guaranteed that bin never exceeds two digits, i.e., 99.
type  arrayUnits is array(0 to 99) of std_logic_vector(3 downto 0);
signal U_Units : arrayUnits := 	("0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001",
			         "0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001",
				 "0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001",
				 "0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001",
				 "0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001",
				 "0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001",
				 "0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001",
				 "0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001",
				 "0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001",
				 "0000", "0001","0010","0011","0100", "0101", "0110", "0111", "1000",  "1001");

type  arrayTens is array(0 to 99) of std_logic_vector(3 downto 0);
signal U_Tens : arrayTens :=  ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000",
			        "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001",
				"0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010", "0010",
				"0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011", "0011",
				"0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100",
				"0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101",
				"0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", 
				"0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", 
				"1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000",
				"1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001");
				
begin
l_bcd<=U_Units(to_integer(unsigned(bin)));
u_bcd <= U_Tens(to_integer(unsigned(bin)));
end architecture rtl;
